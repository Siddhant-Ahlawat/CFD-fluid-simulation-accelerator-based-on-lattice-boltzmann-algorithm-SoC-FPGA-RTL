// Computer_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System (
		input  wire        audio_ADCDAT,                                    //                               audio.ADCDAT
		input  wire        audio_ADCLRCK,                                   //                                    .ADCLRCK
		input  wire        audio_BCLK,                                      //                                    .BCLK
		output wire        audio_DACDAT,                                    //                                    .DACDAT
		input  wire        audio_DACLRCK,                                   //                                    .DACLRCK
		output wire        audio_clk_clk,                                   //                           audio_clk.clk
		input  wire        audio_pll_ref_clk_clk,                           //                   audio_pll_ref_clk.clk
		input  wire        audio_pll_ref_reset_reset,                       //                 audio_pll_ref_reset.reset
		inout  wire        av_config_SDAT,                                  //                           av_config.SDAT
		output wire        av_config_SCLK,                                  //                                    .SCLK
		input  wire [15:0] bus_master_audio_external_interface_address,     // bus_master_audio_external_interface.address
		input  wire [3:0]  bus_master_audio_external_interface_byte_enable, //                                    .byte_enable
		input  wire        bus_master_audio_external_interface_read,        //                                    .read
		input  wire        bus_master_audio_external_interface_write,       //                                    .write
		input  wire [31:0] bus_master_audio_external_interface_write_data,  //                                    .write_data
		output wire        bus_master_audio_external_interface_acknowledge, //                                    .acknowledge
		output wire [31:0] bus_master_audio_external_interface_read_data,   //                                    .read_data
		input  wire [31:0] collide_finish_export,                           //                      collide_finish.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,                 //                              hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,                   //                                    .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,                   //                                    .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,                   //                                    .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,                   //                                    .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,                   //                                    .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,                   //                                    .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,                    //                                    .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,                 //                                    .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,                 //                                    .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,                 //                                    .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,                   //                                    .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,                   //                                    .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,                   //                                    .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,                     //                                    .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,                     //                                    .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,                     //                                    .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,                     //                                    .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,                     //                                    .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,                     //                                    .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                     //                                    .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                      //                                    .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                      //                                    .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,                     //                                    .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                      //                                    .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                      //                                    .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                      //                                    .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                      //                                    .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                      //                                    .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                      //                                    .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                      //                                    .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                      //                                    .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                      //                                    .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                      //                                    .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                     //                                    .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                     //                                    .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                     //                                    .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                     //                                    .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,                    //                                    .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,                   //                                    .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,                   //                                    .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,                    //                                    .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,                     //                                    .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                     //                                    .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,                     //                                    .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,                     //                                    .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,                     //                                    .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,                     //                                    .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,                  //                                    .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,                  //                                    .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,                  //                                    .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,                  //                                    .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,                  //                                    .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,                  //                                    .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,                  //                                    .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,                  //                                    .hps_io_gpio_inst_GPIO61
		input  wire [31:0] init_finish_export,                              //                         init_finish.export
		output wire [31:0] init_ship_export,                                //                           init_ship.export
		output wire [14:0] memory_mem_a,                                    //                              memory.mem_a
		output wire [2:0]  memory_mem_ba,                                   //                                    .mem_ba
		output wire        memory_mem_ck,                                   //                                    .mem_ck
		output wire        memory_mem_ck_n,                                 //                                    .mem_ck_n
		output wire        memory_mem_cke,                                  //                                    .mem_cke
		output wire        memory_mem_cs_n,                                 //                                    .mem_cs_n
		output wire        memory_mem_ras_n,                                //                                    .mem_ras_n
		output wire        memory_mem_cas_n,                                //                                    .mem_cas_n
		output wire        memory_mem_we_n,                                 //                                    .mem_we_n
		output wire        memory_mem_reset_n,                              //                                    .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                   //                                    .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                  //                                    .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                //                                    .mem_dqs_n
		output wire        memory_mem_odt,                                  //                                    .mem_odt
		output wire [3:0]  memory_mem_dm,                                   //                                    .mem_dm
		input  wire        memory_oct_rzqin,                                //                                    .oct_rzqin
		input  wire [31:0] move_trace_finish_export,                        //                   move_trace_finish.export
		output wire [31:0] n0_from_hps_export,                              //                         n0_from_hps.export
		output wire [31:0] ne_from_hps_export,                              //                         ne_from_hps.export
		output wire [31:0] nn_from_hps_export,                              //                         nn_from_hps.export
		output wire [31:0] nne_from_hps_export,                             //                        nne_from_hps.export
		output wire [31:0] nnw_from_hps_export,                             //                        nnw_from_hps.export
		output wire [31:0] ns_from_hps_export,                              //                         ns_from_hps.export
		output wire [31:0] nse_from_hps_export,                             //                        nse_from_hps.export
		output wire [31:0] nsw_from_hps_export,                             //                        nsw_from_hps.export
		output wire [31:0] nw_from_hps_export,                              //                         nw_from_hps.export
		input  wire [31:0] pipes_export,                                    //                               pipes.export
		input  wire [31:0] print_finish_export,                             //                        print_finish.export
		output wire [31:0] reset_lb_export,                                 //                            reset_lb.export
		output wire        sdram_clk_clk,                                   //                           sdram_clk.clk
		output wire [31:0] ship_x_export,                                   //                              ship_x.export
		output wire [31:0] ship_y_export,                                   //                              ship_y.export
		input  wire [31:0] speed_color_finish_export,                       //                  speed_color_finish.export
		output wire [31:0] start_collide_export,                            //                       start_collide.export
		output wire [31:0] start_init_export,                               //                          start_init.export
		output wire [31:0] start_move_trace_export,                         //                    start_move_trace.export
		output wire [31:0] start_print_export,                              //                         start_print.export
		output wire [31:0] start_speed_color_export,                        //                   start_speed_color.export
		output wire [31:0] start_stream_export,                             //                        start_stream.export
		input  wire [31:0] stream_finish_export,                            //                       stream_finish.export
		input  wire        system_pll_ref_clk_clk,                          //                  system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,                      //                system_pll_ref_reset.reset
		output wire [31:0] test_data_export,                                //                           test_data.export
		output wire [31:0] ux_from_hps_export,                              //                         ux_from_hps.export
		input  wire [31:0] ux_in_export,                                    //                               ux_in.export
		output wire [31:0] uy_from_hps_export,                              //                         uy_from_hps.export
		input  wire [31:0] uy_in_export,                                    //                               uy_in.export
		output wire [31:0] write_address_init_export,                       //                  write_address_init.export
		output wire [31:0] x_fish1_export,                                  //                             x_fish1.export
		output wire [31:0] x_fish2_export,                                  //                             x_fish2.export
		output wire [31:0] y_fish1_export,                                  //                             y_fish1.export
		output wire [31:0] y_fish2_export                                   //                             y_fish2.export
	);

	wire         system_pll_sys_clk_clk;                                         // System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, AV_Config:clk, Audio_Subsystem:sys_clk_clk, Bus_master_audio:clk, collide_finish:clk, init_finish:clk, init_ship:clk, mm_interconnect_0:System_PLL_sys_clk_clk, move_trace_finish:clk, n0_from_hps:clk, ne_from_hps:clk, nn_from_hps:clk, nne_from_hps:clk, nnw_from_hps:clk, ns_from_hps:clk, nse_from_hps:clk, nsw_from_hps:clk, nw_from_hps:clk, pipes:clk, print_finish:clk, reset_lb:clk, rst_controller:clk, rst_controller_002:clk, rst_controller_003:clk, ship_x:clk, ship_y:clk, speed_color_finish:clk, start_collide:clk, start_init:clk, start_move_trace:clk, start_print:clk, start_speed_color:clk, start_stream:clk, stream_finish:clk, test_data:clk, ux_from_hps:clk, ux_in:clk, uy_from_hps:clk, uy_in:clk, write_address_init:clk, x_fish1:clk, x_fish2:clk, y_fish1:clk, y_fish2:clk]
	wire  [31:0] bus_master_audio_avalon_master_readdata;                        // mm_interconnect_0:Bus_master_audio_avalon_master_readdata -> Bus_master_audio:avalon_readdata
	wire         bus_master_audio_avalon_master_waitrequest;                     // mm_interconnect_0:Bus_master_audio_avalon_master_waitrequest -> Bus_master_audio:avalon_waitrequest
	wire   [3:0] bus_master_audio_avalon_master_byteenable;                      // Bus_master_audio:avalon_byteenable -> mm_interconnect_0:Bus_master_audio_avalon_master_byteenable
	wire         bus_master_audio_avalon_master_read;                            // Bus_master_audio:avalon_read -> mm_interconnect_0:Bus_master_audio_avalon_master_read
	wire  [15:0] bus_master_audio_avalon_master_address;                         // Bus_master_audio:avalon_address -> mm_interconnect_0:Bus_master_audio_avalon_master_address
	wire         bus_master_audio_avalon_master_write;                           // Bus_master_audio:avalon_write -> mm_interconnect_0:Bus_master_audio_avalon_master_write
	wire  [31:0] bus_master_audio_avalon_master_writedata;                       // Bus_master_audio:avalon_writedata -> mm_interconnect_0:Bus_master_audio_avalon_master_writedata
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                           // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                             // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                             // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire         arm_a9_hps_h2f_lw_axi_master_wready;                            // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                               // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire         arm_a9_hps_h2f_lw_axi_master_rready;                            // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                             // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                               // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                           // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire         arm_a9_hps_h2f_lw_axi_master_wvalid;                            // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                            // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                            // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                            // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                             // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire         arm_a9_hps_h2f_lw_axi_master_arvalid;                           // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                           // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                              // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                            // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                            // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                            // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire         arm_a9_hps_h2f_lw_axi_master_arready;                           // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire         arm_a9_hps_h2f_lw_axi_master_awready;                           // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                           // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                            // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire         arm_a9_hps_h2f_lw_axi_master_bready;                            // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire         arm_a9_hps_h2f_lw_axi_master_rlast;                             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire         arm_a9_hps_h2f_lw_axi_master_wlast;                             // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                              // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                               // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire         arm_a9_hps_h2f_lw_axi_master_bvalid;                            // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                            // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire         arm_a9_hps_h2f_lw_axi_master_awvalid;                           // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire         arm_a9_hps_h2f_lw_axi_master_rvalid;                            // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire         mm_interconnect_0_audio_subsystem_audio_slave_chipselect;       // mm_interconnect_0:Audio_Subsystem_audio_slave_chipselect -> Audio_Subsystem:audio_slave_chipselect
	wire  [31:0] mm_interconnect_0_audio_subsystem_audio_slave_readdata;         // Audio_Subsystem:audio_slave_readdata -> mm_interconnect_0:Audio_Subsystem_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_subsystem_audio_slave_address;          // mm_interconnect_0:Audio_Subsystem_audio_slave_address -> Audio_Subsystem:audio_slave_address
	wire         mm_interconnect_0_audio_subsystem_audio_slave_read;             // mm_interconnect_0:Audio_Subsystem_audio_slave_read -> Audio_Subsystem:audio_slave_read
	wire         mm_interconnect_0_audio_subsystem_audio_slave_write;            // mm_interconnect_0:Audio_Subsystem_audio_slave_write -> Audio_Subsystem:audio_slave_write
	wire  [31:0] mm_interconnect_0_audio_subsystem_audio_slave_writedata;        // mm_interconnect_0:Audio_Subsystem_audio_slave_writedata -> Audio_Subsystem:audio_slave_writedata
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_readdata;    // AV_Config:readdata -> mm_interconnect_0:AV_Config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest; // AV_Config:waitrequest -> mm_interconnect_0:AV_Config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_av_config_avalon_av_config_slave_address;     // mm_interconnect_0:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_read;        // mm_interconnect_0:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	wire   [3:0] mm_interconnect_0_av_config_avalon_av_config_slave_byteenable;  // mm_interconnect_0:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_write;       // mm_interconnect_0:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_writedata;   // mm_interconnect_0:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	wire         mm_interconnect_0_n0_from_hps_s1_chipselect;                    // mm_interconnect_0:n0_from_hps_s1_chipselect -> n0_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_n0_from_hps_s1_readdata;                      // n0_from_hps:readdata -> mm_interconnect_0:n0_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_n0_from_hps_s1_address;                       // mm_interconnect_0:n0_from_hps_s1_address -> n0_from_hps:address
	wire         mm_interconnect_0_n0_from_hps_s1_write;                         // mm_interconnect_0:n0_from_hps_s1_write -> n0_from_hps:write_n
	wire  [31:0] mm_interconnect_0_n0_from_hps_s1_writedata;                     // mm_interconnect_0:n0_from_hps_s1_writedata -> n0_from_hps:writedata
	wire         mm_interconnect_0_nn_from_hps_s1_chipselect;                    // mm_interconnect_0:nn_from_hps_s1_chipselect -> nn_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_nn_from_hps_s1_readdata;                      // nn_from_hps:readdata -> mm_interconnect_0:nn_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_nn_from_hps_s1_address;                       // mm_interconnect_0:nn_from_hps_s1_address -> nn_from_hps:address
	wire         mm_interconnect_0_nn_from_hps_s1_write;                         // mm_interconnect_0:nn_from_hps_s1_write -> nn_from_hps:write_n
	wire  [31:0] mm_interconnect_0_nn_from_hps_s1_writedata;                     // mm_interconnect_0:nn_from_hps_s1_writedata -> nn_from_hps:writedata
	wire         mm_interconnect_0_ns_from_hps_s1_chipselect;                    // mm_interconnect_0:ns_from_hps_s1_chipselect -> ns_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_ns_from_hps_s1_readdata;                      // ns_from_hps:readdata -> mm_interconnect_0:ns_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_ns_from_hps_s1_address;                       // mm_interconnect_0:ns_from_hps_s1_address -> ns_from_hps:address
	wire         mm_interconnect_0_ns_from_hps_s1_write;                         // mm_interconnect_0:ns_from_hps_s1_write -> ns_from_hps:write_n
	wire  [31:0] mm_interconnect_0_ns_from_hps_s1_writedata;                     // mm_interconnect_0:ns_from_hps_s1_writedata -> ns_from_hps:writedata
	wire         mm_interconnect_0_nw_from_hps_s1_chipselect;                    // mm_interconnect_0:nw_from_hps_s1_chipselect -> nw_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_nw_from_hps_s1_readdata;                      // nw_from_hps:readdata -> mm_interconnect_0:nw_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_nw_from_hps_s1_address;                       // mm_interconnect_0:nw_from_hps_s1_address -> nw_from_hps:address
	wire         mm_interconnect_0_nw_from_hps_s1_write;                         // mm_interconnect_0:nw_from_hps_s1_write -> nw_from_hps:write_n
	wire  [31:0] mm_interconnect_0_nw_from_hps_s1_writedata;                     // mm_interconnect_0:nw_from_hps_s1_writedata -> nw_from_hps:writedata
	wire         mm_interconnect_0_ne_from_hps_s1_chipselect;                    // mm_interconnect_0:ne_from_hps_s1_chipselect -> ne_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_ne_from_hps_s1_readdata;                      // ne_from_hps:readdata -> mm_interconnect_0:ne_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_ne_from_hps_s1_address;                       // mm_interconnect_0:ne_from_hps_s1_address -> ne_from_hps:address
	wire         mm_interconnect_0_ne_from_hps_s1_write;                         // mm_interconnect_0:ne_from_hps_s1_write -> ne_from_hps:write_n
	wire  [31:0] mm_interconnect_0_ne_from_hps_s1_writedata;                     // mm_interconnect_0:ne_from_hps_s1_writedata -> ne_from_hps:writedata
	wire         mm_interconnect_0_nnw_from_hps_s1_chipselect;                   // mm_interconnect_0:nnw_from_hps_s1_chipselect -> nnw_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_nnw_from_hps_s1_readdata;                     // nnw_from_hps:readdata -> mm_interconnect_0:nnw_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_nnw_from_hps_s1_address;                      // mm_interconnect_0:nnw_from_hps_s1_address -> nnw_from_hps:address
	wire         mm_interconnect_0_nnw_from_hps_s1_write;                        // mm_interconnect_0:nnw_from_hps_s1_write -> nnw_from_hps:write_n
	wire  [31:0] mm_interconnect_0_nnw_from_hps_s1_writedata;                    // mm_interconnect_0:nnw_from_hps_s1_writedata -> nnw_from_hps:writedata
	wire         mm_interconnect_0_nne_from_hps_s1_chipselect;                   // mm_interconnect_0:nne_from_hps_s1_chipselect -> nne_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_nne_from_hps_s1_readdata;                     // nne_from_hps:readdata -> mm_interconnect_0:nne_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_nne_from_hps_s1_address;                      // mm_interconnect_0:nne_from_hps_s1_address -> nne_from_hps:address
	wire         mm_interconnect_0_nne_from_hps_s1_write;                        // mm_interconnect_0:nne_from_hps_s1_write -> nne_from_hps:write_n
	wire  [31:0] mm_interconnect_0_nne_from_hps_s1_writedata;                    // mm_interconnect_0:nne_from_hps_s1_writedata -> nne_from_hps:writedata
	wire         mm_interconnect_0_nsw_from_hps_s1_chipselect;                   // mm_interconnect_0:nsw_from_hps_s1_chipselect -> nsw_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_nsw_from_hps_s1_readdata;                     // nsw_from_hps:readdata -> mm_interconnect_0:nsw_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_nsw_from_hps_s1_address;                      // mm_interconnect_0:nsw_from_hps_s1_address -> nsw_from_hps:address
	wire         mm_interconnect_0_nsw_from_hps_s1_write;                        // mm_interconnect_0:nsw_from_hps_s1_write -> nsw_from_hps:write_n
	wire  [31:0] mm_interconnect_0_nsw_from_hps_s1_writedata;                    // mm_interconnect_0:nsw_from_hps_s1_writedata -> nsw_from_hps:writedata
	wire         mm_interconnect_0_nse_from_hps_s1_chipselect;                   // mm_interconnect_0:nse_from_hps_s1_chipselect -> nse_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_nse_from_hps_s1_readdata;                     // nse_from_hps:readdata -> mm_interconnect_0:nse_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_nse_from_hps_s1_address;                      // mm_interconnect_0:nse_from_hps_s1_address -> nse_from_hps:address
	wire         mm_interconnect_0_nse_from_hps_s1_write;                        // mm_interconnect_0:nse_from_hps_s1_write -> nse_from_hps:write_n
	wire  [31:0] mm_interconnect_0_nse_from_hps_s1_writedata;                    // mm_interconnect_0:nse_from_hps_s1_writedata -> nse_from_hps:writedata
	wire         mm_interconnect_0_start_collide_s1_chipselect;                  // mm_interconnect_0:start_collide_s1_chipselect -> start_collide:chipselect
	wire  [31:0] mm_interconnect_0_start_collide_s1_readdata;                    // start_collide:readdata -> mm_interconnect_0:start_collide_s1_readdata
	wire   [1:0] mm_interconnect_0_start_collide_s1_address;                     // mm_interconnect_0:start_collide_s1_address -> start_collide:address
	wire         mm_interconnect_0_start_collide_s1_write;                       // mm_interconnect_0:start_collide_s1_write -> start_collide:write_n
	wire  [31:0] mm_interconnect_0_start_collide_s1_writedata;                   // mm_interconnect_0:start_collide_s1_writedata -> start_collide:writedata
	wire  [31:0] mm_interconnect_0_collide_finish_s1_readdata;                   // collide_finish:readdata -> mm_interconnect_0:collide_finish_s1_readdata
	wire   [1:0] mm_interconnect_0_collide_finish_s1_address;                    // mm_interconnect_0:collide_finish_s1_address -> collide_finish:address
	wire         mm_interconnect_0_start_stream_s1_chipselect;                   // mm_interconnect_0:start_stream_s1_chipselect -> start_stream:chipselect
	wire  [31:0] mm_interconnect_0_start_stream_s1_readdata;                     // start_stream:readdata -> mm_interconnect_0:start_stream_s1_readdata
	wire   [1:0] mm_interconnect_0_start_stream_s1_address;                      // mm_interconnect_0:start_stream_s1_address -> start_stream:address
	wire         mm_interconnect_0_start_stream_s1_write;                        // mm_interconnect_0:start_stream_s1_write -> start_stream:write_n
	wire  [31:0] mm_interconnect_0_start_stream_s1_writedata;                    // mm_interconnect_0:start_stream_s1_writedata -> start_stream:writedata
	wire  [31:0] mm_interconnect_0_stream_finish_s1_readdata;                    // stream_finish:readdata -> mm_interconnect_0:stream_finish_s1_readdata
	wire   [1:0] mm_interconnect_0_stream_finish_s1_address;                     // mm_interconnect_0:stream_finish_s1_address -> stream_finish:address
	wire         mm_interconnect_0_write_address_init_s1_chipselect;             // mm_interconnect_0:write_address_init_s1_chipselect -> write_address_init:chipselect
	wire  [31:0] mm_interconnect_0_write_address_init_s1_readdata;               // write_address_init:readdata -> mm_interconnect_0:write_address_init_s1_readdata
	wire   [1:0] mm_interconnect_0_write_address_init_s1_address;                // mm_interconnect_0:write_address_init_s1_address -> write_address_init:address
	wire         mm_interconnect_0_write_address_init_s1_write;                  // mm_interconnect_0:write_address_init_s1_write -> write_address_init:write_n
	wire  [31:0] mm_interconnect_0_write_address_init_s1_writedata;              // mm_interconnect_0:write_address_init_s1_writedata -> write_address_init:writedata
	wire         mm_interconnect_0_start_init_s1_chipselect;                     // mm_interconnect_0:start_init_s1_chipselect -> start_init:chipselect
	wire  [31:0] mm_interconnect_0_start_init_s1_readdata;                       // start_init:readdata -> mm_interconnect_0:start_init_s1_readdata
	wire   [1:0] mm_interconnect_0_start_init_s1_address;                        // mm_interconnect_0:start_init_s1_address -> start_init:address
	wire         mm_interconnect_0_start_init_s1_write;                          // mm_interconnect_0:start_init_s1_write -> start_init:write_n
	wire  [31:0] mm_interconnect_0_start_init_s1_writedata;                      // mm_interconnect_0:start_init_s1_writedata -> start_init:writedata
	wire  [31:0] mm_interconnect_0_init_finish_s1_readdata;                      // init_finish:readdata -> mm_interconnect_0:init_finish_s1_readdata
	wire   [1:0] mm_interconnect_0_init_finish_s1_address;                       // mm_interconnect_0:init_finish_s1_address -> init_finish:address
	wire         mm_interconnect_0_init_ship_s1_chipselect;                      // mm_interconnect_0:init_ship_s1_chipselect -> init_ship:chipselect
	wire  [31:0] mm_interconnect_0_init_ship_s1_readdata;                        // init_ship:readdata -> mm_interconnect_0:init_ship_s1_readdata
	wire   [1:0] mm_interconnect_0_init_ship_s1_address;                         // mm_interconnect_0:init_ship_s1_address -> init_ship:address
	wire         mm_interconnect_0_init_ship_s1_write;                           // mm_interconnect_0:init_ship_s1_write -> init_ship:write_n
	wire  [31:0] mm_interconnect_0_init_ship_s1_writedata;                       // mm_interconnect_0:init_ship_s1_writedata -> init_ship:writedata
	wire         mm_interconnect_0_start_move_trace_s1_chipselect;               // mm_interconnect_0:start_move_trace_s1_chipselect -> start_move_trace:chipselect
	wire  [31:0] mm_interconnect_0_start_move_trace_s1_readdata;                 // start_move_trace:readdata -> mm_interconnect_0:start_move_trace_s1_readdata
	wire   [1:0] mm_interconnect_0_start_move_trace_s1_address;                  // mm_interconnect_0:start_move_trace_s1_address -> start_move_trace:address
	wire         mm_interconnect_0_start_move_trace_s1_write;                    // mm_interconnect_0:start_move_trace_s1_write -> start_move_trace:write_n
	wire  [31:0] mm_interconnect_0_start_move_trace_s1_writedata;                // mm_interconnect_0:start_move_trace_s1_writedata -> start_move_trace:writedata
	wire  [31:0] mm_interconnect_0_move_trace_finish_s1_readdata;                // move_trace_finish:readdata -> mm_interconnect_0:move_trace_finish_s1_readdata
	wire   [1:0] mm_interconnect_0_move_trace_finish_s1_address;                 // mm_interconnect_0:move_trace_finish_s1_address -> move_trace_finish:address
	wire         mm_interconnect_0_start_speed_color_s1_chipselect;              // mm_interconnect_0:start_speed_color_s1_chipselect -> start_speed_color:chipselect
	wire  [31:0] mm_interconnect_0_start_speed_color_s1_readdata;                // start_speed_color:readdata -> mm_interconnect_0:start_speed_color_s1_readdata
	wire   [1:0] mm_interconnect_0_start_speed_color_s1_address;                 // mm_interconnect_0:start_speed_color_s1_address -> start_speed_color:address
	wire         mm_interconnect_0_start_speed_color_s1_write;                   // mm_interconnect_0:start_speed_color_s1_write -> start_speed_color:write_n
	wire  [31:0] mm_interconnect_0_start_speed_color_s1_writedata;               // mm_interconnect_0:start_speed_color_s1_writedata -> start_speed_color:writedata
	wire  [31:0] mm_interconnect_0_speed_color_finish_s1_readdata;               // speed_color_finish:readdata -> mm_interconnect_0:speed_color_finish_s1_readdata
	wire   [1:0] mm_interconnect_0_speed_color_finish_s1_address;                // mm_interconnect_0:speed_color_finish_s1_address -> speed_color_finish:address
	wire         mm_interconnect_0_ux_from_hps_s1_chipselect;                    // mm_interconnect_0:ux_from_hps_s1_chipselect -> ux_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_ux_from_hps_s1_readdata;                      // ux_from_hps:readdata -> mm_interconnect_0:ux_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_ux_from_hps_s1_address;                       // mm_interconnect_0:ux_from_hps_s1_address -> ux_from_hps:address
	wire         mm_interconnect_0_ux_from_hps_s1_write;                         // mm_interconnect_0:ux_from_hps_s1_write -> ux_from_hps:write_n
	wire  [31:0] mm_interconnect_0_ux_from_hps_s1_writedata;                     // mm_interconnect_0:ux_from_hps_s1_writedata -> ux_from_hps:writedata
	wire         mm_interconnect_0_uy_from_hps_s1_chipselect;                    // mm_interconnect_0:uy_from_hps_s1_chipselect -> uy_from_hps:chipselect
	wire  [31:0] mm_interconnect_0_uy_from_hps_s1_readdata;                      // uy_from_hps:readdata -> mm_interconnect_0:uy_from_hps_s1_readdata
	wire   [1:0] mm_interconnect_0_uy_from_hps_s1_address;                       // mm_interconnect_0:uy_from_hps_s1_address -> uy_from_hps:address
	wire         mm_interconnect_0_uy_from_hps_s1_write;                         // mm_interconnect_0:uy_from_hps_s1_write -> uy_from_hps:write_n
	wire  [31:0] mm_interconnect_0_uy_from_hps_s1_writedata;                     // mm_interconnect_0:uy_from_hps_s1_writedata -> uy_from_hps:writedata
	wire         mm_interconnect_0_reset_lb_s1_chipselect;                       // mm_interconnect_0:reset_lb_s1_chipselect -> reset_lb:chipselect
	wire  [31:0] mm_interconnect_0_reset_lb_s1_readdata;                         // reset_lb:readdata -> mm_interconnect_0:reset_lb_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_lb_s1_address;                          // mm_interconnect_0:reset_lb_s1_address -> reset_lb:address
	wire         mm_interconnect_0_reset_lb_s1_write;                            // mm_interconnect_0:reset_lb_s1_write -> reset_lb:write_n
	wire  [31:0] mm_interconnect_0_reset_lb_s1_writedata;                        // mm_interconnect_0:reset_lb_s1_writedata -> reset_lb:writedata
	wire  [31:0] mm_interconnect_0_pipes_s1_readdata;                            // pipes:readdata -> mm_interconnect_0:pipes_s1_readdata
	wire   [1:0] mm_interconnect_0_pipes_s1_address;                             // mm_interconnect_0:pipes_s1_address -> pipes:address
	wire         mm_interconnect_0_start_print_s1_chipselect;                    // mm_interconnect_0:start_print_s1_chipselect -> start_print:chipselect
	wire  [31:0] mm_interconnect_0_start_print_s1_readdata;                      // start_print:readdata -> mm_interconnect_0:start_print_s1_readdata
	wire   [1:0] mm_interconnect_0_start_print_s1_address;                       // mm_interconnect_0:start_print_s1_address -> start_print:address
	wire         mm_interconnect_0_start_print_s1_write;                         // mm_interconnect_0:start_print_s1_write -> start_print:write_n
	wire  [31:0] mm_interconnect_0_start_print_s1_writedata;                     // mm_interconnect_0:start_print_s1_writedata -> start_print:writedata
	wire  [31:0] mm_interconnect_0_print_finish_s1_readdata;                     // print_finish:readdata -> mm_interconnect_0:print_finish_s1_readdata
	wire   [1:0] mm_interconnect_0_print_finish_s1_address;                      // mm_interconnect_0:print_finish_s1_address -> print_finish:address
	wire         mm_interconnect_0_test_data_s1_chipselect;                      // mm_interconnect_0:test_data_s1_chipselect -> test_data:chipselect
	wire  [31:0] mm_interconnect_0_test_data_s1_readdata;                        // test_data:readdata -> mm_interconnect_0:test_data_s1_readdata
	wire   [1:0] mm_interconnect_0_test_data_s1_address;                         // mm_interconnect_0:test_data_s1_address -> test_data:address
	wire         mm_interconnect_0_test_data_s1_write;                           // mm_interconnect_0:test_data_s1_write -> test_data:write_n
	wire  [31:0] mm_interconnect_0_test_data_s1_writedata;                       // mm_interconnect_0:test_data_s1_writedata -> test_data:writedata
	wire         mm_interconnect_0_ship_x_s1_chipselect;                         // mm_interconnect_0:ship_x_s1_chipselect -> ship_x:chipselect
	wire  [31:0] mm_interconnect_0_ship_x_s1_readdata;                           // ship_x:readdata -> mm_interconnect_0:ship_x_s1_readdata
	wire   [1:0] mm_interconnect_0_ship_x_s1_address;                            // mm_interconnect_0:ship_x_s1_address -> ship_x:address
	wire         mm_interconnect_0_ship_x_s1_write;                              // mm_interconnect_0:ship_x_s1_write -> ship_x:write_n
	wire  [31:0] mm_interconnect_0_ship_x_s1_writedata;                          // mm_interconnect_0:ship_x_s1_writedata -> ship_x:writedata
	wire         mm_interconnect_0_ship_y_s1_chipselect;                         // mm_interconnect_0:ship_y_s1_chipselect -> ship_y:chipselect
	wire  [31:0] mm_interconnect_0_ship_y_s1_readdata;                           // ship_y:readdata -> mm_interconnect_0:ship_y_s1_readdata
	wire   [1:0] mm_interconnect_0_ship_y_s1_address;                            // mm_interconnect_0:ship_y_s1_address -> ship_y:address
	wire         mm_interconnect_0_ship_y_s1_write;                              // mm_interconnect_0:ship_y_s1_write -> ship_y:write_n
	wire  [31:0] mm_interconnect_0_ship_y_s1_writedata;                          // mm_interconnect_0:ship_y_s1_writedata -> ship_y:writedata
	wire  [31:0] mm_interconnect_0_ux_in_s1_readdata;                            // ux_in:readdata -> mm_interconnect_0:ux_in_s1_readdata
	wire   [1:0] mm_interconnect_0_ux_in_s1_address;                             // mm_interconnect_0:ux_in_s1_address -> ux_in:address
	wire  [31:0] mm_interconnect_0_uy_in_s1_readdata;                            // uy_in:readdata -> mm_interconnect_0:uy_in_s1_readdata
	wire   [1:0] mm_interconnect_0_uy_in_s1_address;                             // mm_interconnect_0:uy_in_s1_address -> uy_in:address
	wire         mm_interconnect_0_x_fish1_s1_chipselect;                        // mm_interconnect_0:x_fish1_s1_chipselect -> x_fish1:chipselect
	wire  [31:0] mm_interconnect_0_x_fish1_s1_readdata;                          // x_fish1:readdata -> mm_interconnect_0:x_fish1_s1_readdata
	wire   [1:0] mm_interconnect_0_x_fish1_s1_address;                           // mm_interconnect_0:x_fish1_s1_address -> x_fish1:address
	wire         mm_interconnect_0_x_fish1_s1_write;                             // mm_interconnect_0:x_fish1_s1_write -> x_fish1:write_n
	wire  [31:0] mm_interconnect_0_x_fish1_s1_writedata;                         // mm_interconnect_0:x_fish1_s1_writedata -> x_fish1:writedata
	wire         mm_interconnect_0_y_fish1_s1_chipselect;                        // mm_interconnect_0:y_fish1_s1_chipselect -> y_fish1:chipselect
	wire  [31:0] mm_interconnect_0_y_fish1_s1_readdata;                          // y_fish1:readdata -> mm_interconnect_0:y_fish1_s1_readdata
	wire   [1:0] mm_interconnect_0_y_fish1_s1_address;                           // mm_interconnect_0:y_fish1_s1_address -> y_fish1:address
	wire         mm_interconnect_0_y_fish1_s1_write;                             // mm_interconnect_0:y_fish1_s1_write -> y_fish1:write_n
	wire  [31:0] mm_interconnect_0_y_fish1_s1_writedata;                         // mm_interconnect_0:y_fish1_s1_writedata -> y_fish1:writedata
	wire         mm_interconnect_0_x_fish2_s1_chipselect;                        // mm_interconnect_0:x_fish2_s1_chipselect -> x_fish2:chipselect
	wire  [31:0] mm_interconnect_0_x_fish2_s1_readdata;                          // x_fish2:readdata -> mm_interconnect_0:x_fish2_s1_readdata
	wire   [1:0] mm_interconnect_0_x_fish2_s1_address;                           // mm_interconnect_0:x_fish2_s1_address -> x_fish2:address
	wire         mm_interconnect_0_x_fish2_s1_write;                             // mm_interconnect_0:x_fish2_s1_write -> x_fish2:write_n
	wire  [31:0] mm_interconnect_0_x_fish2_s1_writedata;                         // mm_interconnect_0:x_fish2_s1_writedata -> x_fish2:writedata
	wire         mm_interconnect_0_y_fish2_s1_chipselect;                        // mm_interconnect_0:y_fish2_s1_chipselect -> y_fish2:chipselect
	wire  [31:0] mm_interconnect_0_y_fish2_s1_readdata;                          // y_fish2:readdata -> mm_interconnect_0:y_fish2_s1_readdata
	wire   [1:0] mm_interconnect_0_y_fish2_s1_address;                           // mm_interconnect_0:y_fish2_s1_address -> y_fish2:address
	wire         mm_interconnect_0_y_fish2_s1_write;                             // mm_interconnect_0:y_fish2_s1_write -> y_fish2:write_n
	wire  [31:0] mm_interconnect_0_y_fish2_s1_writedata;                         // mm_interconnect_0:y_fish2_s1_writedata -> y_fish2:writedata
	wire         irq_mapper_receiver0_irq;                                       // Audio_Subsystem:audio_irq_irq -> irq_mapper:receiver0_irq
	wire  [31:0] arm_a9_hps_f2h_irq0_irq;                                        // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;                                        // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [AV_Config:reset, Bus_master_audio:reset, mm_interconnect_0:Audio_Subsystem_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_0:Bus_master_audio_reset_reset_bridge_in_reset_reset]
	wire         arm_a9_hps_h2f_reset_reset;                                     // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_003:reset_in0]
	wire         system_pll_reset_source_reset;                                  // System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> Audio_Subsystem:sys_reset_reset_n
	wire         rst_controller_002_reset_out_reset;                             // rst_controller_002:reset_out -> [collide_finish:reset_n, init_finish:reset_n, init_ship:reset_n, mm_interconnect_0:n0_from_hps_reset_reset_bridge_in_reset_reset, move_trace_finish:reset_n, n0_from_hps:reset_n, ne_from_hps:reset_n, nn_from_hps:reset_n, nne_from_hps:reset_n, nnw_from_hps:reset_n, ns_from_hps:reset_n, nse_from_hps:reset_n, nsw_from_hps:reset_n, nw_from_hps:reset_n, pipes:reset_n, print_finish:reset_n, reset_lb:reset_n, ship_x:reset_n, ship_y:reset_n, speed_color_finish:reset_n, start_collide:reset_n, start_init:reset_n, start_move_trace:reset_n, start_print:reset_n, start_speed_color:reset_n, start_stream:reset_n, stream_finish:reset_n, test_data:reset_n, ux_from_hps:reset_n, ux_in:reset_n, uy_from_hps:reset_n, uy_in:reset_n, write_address_init:reset_n, x_fish1:reset_n, x_fish2:reset_n, y_fish1:reset_n, y_fish2:reset_n]
	wire         rst_controller_003_reset_out_reset;                             // rst_controller_003:reset_out -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                         //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                        //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                        //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                      //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                       //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                      //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                     //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                     //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                      //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                   //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                        //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                       //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                     //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                       //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                        //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                     //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),      //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),        //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),        //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),        //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),        //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),        //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),        //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),         //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),      //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),      //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),      //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),        //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),        //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),        //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),          //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),          //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),          //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),          //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),          //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),          //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),          //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),           //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),           //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),          //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),           //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),           //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),           //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),           //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),           //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),           //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),           //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),           //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),           //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),           //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),          //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),          //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),          //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),          //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),         //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),        //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),        //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),         //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),          //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),          //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),          //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),          //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),          //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),          //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),       //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),       //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),       //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),       //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),       //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),       //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),       //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),       //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),               //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                     //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                     //                  .awaddr
		.h2f_AWLEN                (),                                     //                  .awlen
		.h2f_AWSIZE               (),                                     //                  .awsize
		.h2f_AWBURST              (),                                     //                  .awburst
		.h2f_AWLOCK               (),                                     //                  .awlock
		.h2f_AWCACHE              (),                                     //                  .awcache
		.h2f_AWPROT               (),                                     //                  .awprot
		.h2f_AWVALID              (),                                     //                  .awvalid
		.h2f_AWREADY              (),                                     //                  .awready
		.h2f_WID                  (),                                     //                  .wid
		.h2f_WDATA                (),                                     //                  .wdata
		.h2f_WSTRB                (),                                     //                  .wstrb
		.h2f_WLAST                (),                                     //                  .wlast
		.h2f_WVALID               (),                                     //                  .wvalid
		.h2f_WREADY               (),                                     //                  .wready
		.h2f_BID                  (),                                     //                  .bid
		.h2f_BRESP                (),                                     //                  .bresp
		.h2f_BVALID               (),                                     //                  .bvalid
		.h2f_BREADY               (),                                     //                  .bready
		.h2f_ARID                 (),                                     //                  .arid
		.h2f_ARADDR               (),                                     //                  .araddr
		.h2f_ARLEN                (),                                     //                  .arlen
		.h2f_ARSIZE               (),                                     //                  .arsize
		.h2f_ARBURST              (),                                     //                  .arburst
		.h2f_ARLOCK               (),                                     //                  .arlock
		.h2f_ARCACHE              (),                                     //                  .arcache
		.h2f_ARPROT               (),                                     //                  .arprot
		.h2f_ARVALID              (),                                     //                  .arvalid
		.h2f_ARREADY              (),                                     //                  .arready
		.h2f_RID                  (),                                     //                  .rid
		.h2f_RDATA                (),                                     //                  .rdata
		.h2f_RRESP                (),                                     //                  .rresp
		.h2f_RLAST                (),                                     //                  .rlast
		.h2f_RVALID               (),                                     //                  .rvalid
		.h2f_RREADY               (),                                     //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),               //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                     //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                     //                  .awaddr
		.f2h_AWLEN                (),                                     //                  .awlen
		.f2h_AWSIZE               (),                                     //                  .awsize
		.f2h_AWBURST              (),                                     //                  .awburst
		.f2h_AWLOCK               (),                                     //                  .awlock
		.f2h_AWCACHE              (),                                     //                  .awcache
		.f2h_AWPROT               (),                                     //                  .awprot
		.f2h_AWVALID              (),                                     //                  .awvalid
		.f2h_AWREADY              (),                                     //                  .awready
		.f2h_AWUSER               (),                                     //                  .awuser
		.f2h_WID                  (),                                     //                  .wid
		.f2h_WDATA                (),                                     //                  .wdata
		.f2h_WSTRB                (),                                     //                  .wstrb
		.f2h_WLAST                (),                                     //                  .wlast
		.f2h_WVALID               (),                                     //                  .wvalid
		.f2h_WREADY               (),                                     //                  .wready
		.f2h_BID                  (),                                     //                  .bid
		.f2h_BRESP                (),                                     //                  .bresp
		.f2h_BVALID               (),                                     //                  .bvalid
		.f2h_BREADY               (),                                     //                  .bready
		.f2h_ARID                 (),                                     //                  .arid
		.f2h_ARADDR               (),                                     //                  .araddr
		.f2h_ARLEN                (),                                     //                  .arlen
		.f2h_ARSIZE               (),                                     //                  .arsize
		.f2h_ARBURST              (),                                     //                  .arburst
		.f2h_ARLOCK               (),                                     //                  .arlock
		.f2h_ARCACHE              (),                                     //                  .arcache
		.f2h_ARPROT               (),                                     //                  .arprot
		.f2h_ARVALID              (),                                     //                  .arvalid
		.f2h_ARREADY              (),                                     //                  .arready
		.f2h_ARUSER               (),                                     //                  .aruser
		.f2h_RID                  (),                                     //                  .rid
		.f2h_RDATA                (),                                     //                  .rdata
		.f2h_RRESP                (),                                     //                  .rresp
		.f2h_RLAST                (),                                     //                  .rlast
		.f2h_RVALID               (),                                     //                  .rvalid
		.f2h_RREADY               (),                                     //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	Computer_System_AV_Config av_config (
		.clk         (system_pll_sys_clk_clk),                                         //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //                  reset.reset
		.address     (mm_interconnect_0_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (av_config_SDAT),                                                 //     external_interface.export
		.I2C_SCLK    (av_config_SCLK)                                                  //                       .export
	);

	Computer_System_Audio_Subsystem audio_subsystem (
		.audio_ADCDAT              (audio_ADCDAT),                                             //               audio.ADCDAT
		.audio_ADCLRCK             (audio_ADCLRCK),                                            //                    .ADCLRCK
		.audio_BCLK                (audio_BCLK),                                               //                    .BCLK
		.audio_DACDAT              (audio_DACDAT),                                             //                    .DACDAT
		.audio_DACLRCK             (audio_DACLRCK),                                            //                    .DACLRCK
		.audio_clk_clk             (audio_clk_clk),                                            //           audio_clk.clk
		.audio_irq_irq             (irq_mapper_receiver0_irq),                                 //           audio_irq.irq
		.audio_pll_ref_clk_clk     (audio_pll_ref_clk_clk),                                    //   audio_pll_ref_clk.clk
		.audio_pll_ref_reset_reset (audio_pll_ref_reset_reset),                                // audio_pll_ref_reset.reset
		.audio_reset_reset         (),                                                         //         audio_reset.reset
		.audio_slave_address       (mm_interconnect_0_audio_subsystem_audio_slave_address),    //         audio_slave.address
		.audio_slave_chipselect    (mm_interconnect_0_audio_subsystem_audio_slave_chipselect), //                    .chipselect
		.audio_slave_read          (mm_interconnect_0_audio_subsystem_audio_slave_read),       //                    .read
		.audio_slave_write         (mm_interconnect_0_audio_subsystem_audio_slave_write),      //                    .write
		.audio_slave_writedata     (mm_interconnect_0_audio_subsystem_audio_slave_writedata),  //                    .writedata
		.audio_slave_readdata      (mm_interconnect_0_audio_subsystem_audio_slave_readdata),   //                    .readdata
		.sys_clk_clk               (system_pll_sys_clk_clk),                                   //             sys_clk.clk
		.sys_reset_reset_n         (~rst_controller_001_reset_out_reset)                       //           sys_reset.reset_n
	);

	Computer_System_Bus_master_audio bus_master_audio (
		.clk                (system_pll_sys_clk_clk),                          //                clk.clk
		.reset              (rst_controller_reset_out_reset),                  //              reset.reset
		.avalon_readdata    (bus_master_audio_avalon_master_readdata),         //      avalon_master.readdata
		.avalon_waitrequest (bus_master_audio_avalon_master_waitrequest),      //                   .waitrequest
		.avalon_byteenable  (bus_master_audio_avalon_master_byteenable),       //                   .byteenable
		.avalon_read        (bus_master_audio_avalon_master_read),             //                   .read
		.avalon_write       (bus_master_audio_avalon_master_write),            //                   .write
		.avalon_writedata   (bus_master_audio_avalon_master_writedata),        //                   .writedata
		.avalon_address     (bus_master_audio_avalon_master_address),          //                   .address
		.address            (bus_master_audio_external_interface_address),     // external_interface.export
		.byte_enable        (bus_master_audio_external_interface_byte_enable), //                   .export
		.read               (bus_master_audio_external_interface_read),        //                   .export
		.write              (bus_master_audio_external_interface_write),       //                   .export
		.write_data         (bus_master_audio_external_interface_write_data),  //                   .export
		.acknowledge        (bus_master_audio_external_interface_acknowledge), //                   .export
		.read_data          (bus_master_audio_external_interface_read_data)    //                   .export
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_collide_finish collide_finish (
		.clk      (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_collide_finish_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_collide_finish_s1_readdata), //                    .readdata
		.in_port  (collide_finish_export)                         // external_connection.export
	);

	Computer_System_collide_finish init_finish (
		.clk      (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_init_finish_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_init_finish_s1_readdata), //                    .readdata
		.in_port  (init_finish_export)                         // external_connection.export
	);

	Computer_System_init_ship init_ship (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_init_ship_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_init_ship_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_init_ship_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_init_ship_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_init_ship_s1_readdata),   //                    .readdata
		.out_port   (init_ship_export)                           // external_connection.export
	);

	Computer_System_collide_finish move_trace_finish (
		.clk      (system_pll_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_move_trace_finish_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_move_trace_finish_s1_readdata), //                    .readdata
		.in_port  (move_trace_finish_export)                         // external_connection.export
	);

	Computer_System_init_ship n0_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_n0_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_n0_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_n0_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_n0_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_n0_from_hps_s1_readdata),   //                    .readdata
		.out_port   (n0_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship ne_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_ne_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ne_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ne_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ne_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ne_from_hps_s1_readdata),   //                    .readdata
		.out_port   (ne_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship nn_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_nn_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nn_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nn_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nn_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nn_from_hps_s1_readdata),   //                    .readdata
		.out_port   (nn_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship nne_from_hps (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_nne_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nne_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nne_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nne_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nne_from_hps_s1_readdata),   //                    .readdata
		.out_port   (nne_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship nnw_from_hps (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_nnw_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nnw_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nnw_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nnw_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nnw_from_hps_s1_readdata),   //                    .readdata
		.out_port   (nnw_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship ns_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_ns_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ns_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ns_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ns_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ns_from_hps_s1_readdata),   //                    .readdata
		.out_port   (ns_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship nse_from_hps (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_nse_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nse_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nse_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nse_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nse_from_hps_s1_readdata),   //                    .readdata
		.out_port   (nse_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship nsw_from_hps (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_nsw_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nsw_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nsw_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nsw_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nsw_from_hps_s1_readdata),   //                    .readdata
		.out_port   (nsw_from_hps_export)                           // external_connection.export
	);

	Computer_System_init_ship nw_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_nw_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nw_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nw_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nw_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nw_from_hps_s1_readdata),   //                    .readdata
		.out_port   (nw_from_hps_export)                           // external_connection.export
	);

	Computer_System_collide_finish pipes (
		.clk      (system_pll_sys_clk_clk),              //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_pipes_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pipes_s1_readdata), //                    .readdata
		.in_port  (pipes_export)                         // external_connection.export
	);

	Computer_System_collide_finish print_finish (
		.clk      (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_print_finish_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_print_finish_s1_readdata), //                    .readdata
		.in_port  (print_finish_export)                         // external_connection.export
	);

	Computer_System_init_ship reset_lb (
		.clk        (system_pll_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_reset_lb_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_lb_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_lb_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_lb_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_lb_s1_readdata),   //                    .readdata
		.out_port   (reset_lb_export)                           // external_connection.export
	);

	Computer_System_init_ship ship_x (
		.clk        (system_pll_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_ship_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ship_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ship_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ship_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ship_x_s1_readdata),   //                    .readdata
		.out_port   (ship_x_export)                           // external_connection.export
	);

	Computer_System_init_ship ship_y (
		.clk        (system_pll_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_ship_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ship_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ship_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ship_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ship_y_s1_readdata),   //                    .readdata
		.out_port   (ship_y_export)                           // external_connection.export
	);

	Computer_System_collide_finish speed_color_finish (
		.clk      (system_pll_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_speed_color_finish_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_speed_color_finish_s1_readdata), //                    .readdata
		.in_port  (speed_color_finish_export)                         // external_connection.export
	);

	Computer_System_init_ship start_collide (
		.clk        (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_start_collide_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_collide_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_collide_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_collide_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_collide_s1_readdata),   //                    .readdata
		.out_port   (start_collide_export)                           // external_connection.export
	);

	Computer_System_init_ship start_init (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_start_init_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_init_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_init_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_init_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_init_s1_readdata),   //                    .readdata
		.out_port   (start_init_export)                           // external_connection.export
	);

	Computer_System_init_ship start_move_trace (
		.clk        (system_pll_sys_clk_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_start_move_trace_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_move_trace_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_move_trace_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_move_trace_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_move_trace_s1_readdata),   //                    .readdata
		.out_port   (start_move_trace_export)                           // external_connection.export
	);

	Computer_System_init_ship start_print (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_start_print_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_print_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_print_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_print_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_print_s1_readdata),   //                    .readdata
		.out_port   (start_print_export)                           // external_connection.export
	);

	Computer_System_init_ship start_speed_color (
		.clk        (system_pll_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_start_speed_color_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_speed_color_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_speed_color_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_speed_color_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_speed_color_s1_readdata),   //                    .readdata
		.out_port   (start_speed_color_export)                           // external_connection.export
	);

	Computer_System_init_ship start_stream (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_start_stream_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_stream_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_stream_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_stream_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_stream_s1_readdata),   //                    .readdata
		.out_port   (start_stream_export)                           // external_connection.export
	);

	Computer_System_collide_finish stream_finish (
		.clk      (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_stream_finish_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_stream_finish_s1_readdata), //                    .readdata
		.in_port  (stream_finish_export)                         // external_connection.export
	);

	Computer_System_init_ship test_data (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_test_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_test_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_test_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_test_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_test_data_s1_readdata),   //                    .readdata
		.out_port   (test_data_export)                           // external_connection.export
	);

	Computer_System_init_ship ux_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_ux_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ux_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ux_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ux_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ux_from_hps_s1_readdata),   //                    .readdata
		.out_port   (ux_from_hps_export)                           // external_connection.export
	);

	Computer_System_collide_finish ux_in (
		.clk      (system_pll_sys_clk_clk),              //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_ux_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ux_in_s1_readdata), //                    .readdata
		.in_port  (ux_in_export)                         // external_connection.export
	);

	Computer_System_init_ship uy_from_hps (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_uy_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_uy_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_uy_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_uy_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_uy_from_hps_s1_readdata),   //                    .readdata
		.out_port   (uy_from_hps_export)                           // external_connection.export
	);

	Computer_System_collide_finish uy_in (
		.clk      (system_pll_sys_clk_clk),              //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_uy_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_uy_in_s1_readdata), //                    .readdata
		.in_port  (uy_in_export)                         // external_connection.export
	);

	Computer_System_init_ship write_address_init (
		.clk        (system_pll_sys_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_write_address_init_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_write_address_init_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_write_address_init_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_write_address_init_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_write_address_init_s1_readdata),   //                    .readdata
		.out_port   (write_address_init_export)                           // external_connection.export
	);

	Computer_System_init_ship x_fish1 (
		.clk        (system_pll_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_x_fish1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_x_fish1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_x_fish1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_x_fish1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_x_fish1_s1_readdata),   //                    .readdata
		.out_port   (x_fish1_export)                           // external_connection.export
	);

	Computer_System_init_ship x_fish2 (
		.clk        (system_pll_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_x_fish2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_x_fish2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_x_fish2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_x_fish2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_x_fish2_s1_readdata),   //                    .readdata
		.out_port   (x_fish2_export)                           // external_connection.export
	);

	Computer_System_init_ship y_fish1 (
		.clk        (system_pll_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_y_fish1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_y_fish1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_y_fish1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_y_fish1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_y_fish1_s1_readdata),   //                    .readdata
		.out_port   (y_fish1_export)                           // external_connection.export
	);

	Computer_System_init_ship y_fish2 (
		.clk        (system_pll_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_y_fish2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_y_fish2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_y_fish2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_y_fish2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_y_fish2_s1_readdata),   //                    .readdata
		.out_port   (y_fish2_export)                           // external_connection.export
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                              //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                            //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                             //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                            //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                           //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                            //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                           //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                            //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                           //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                           //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                               //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                             //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                             //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                             //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                            //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                            //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                               //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                             //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                            //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                            //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                              //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                            //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                             //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                            //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                           //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                            //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                           //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                            //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                           //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                           //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                               //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                             //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                             //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                             //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                            //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                            //                                                                   .rready
		.System_PLL_sys_clk_clk                                                   (system_pll_sys_clk_clk),                                         //                                                 System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                             // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Audio_Subsystem_sys_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                                 //                    Audio_Subsystem_sys_reset_reset_bridge_in_reset.reset
		.Bus_master_audio_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                                 //                       Bus_master_audio_reset_reset_bridge_in_reset.reset
		.n0_from_hps_reset_reset_bridge_in_reset_reset                            (rst_controller_002_reset_out_reset),                             //                            n0_from_hps_reset_reset_bridge_in_reset.reset
		.Bus_master_audio_avalon_master_address                                   (bus_master_audio_avalon_master_address),                         //                                     Bus_master_audio_avalon_master.address
		.Bus_master_audio_avalon_master_waitrequest                               (bus_master_audio_avalon_master_waitrequest),                     //                                                                   .waitrequest
		.Bus_master_audio_avalon_master_byteenable                                (bus_master_audio_avalon_master_byteenable),                      //                                                                   .byteenable
		.Bus_master_audio_avalon_master_read                                      (bus_master_audio_avalon_master_read),                            //                                                                   .read
		.Bus_master_audio_avalon_master_readdata                                  (bus_master_audio_avalon_master_readdata),                        //                                                                   .readdata
		.Bus_master_audio_avalon_master_write                                     (bus_master_audio_avalon_master_write),                           //                                                                   .write
		.Bus_master_audio_avalon_master_writedata                                 (bus_master_audio_avalon_master_writedata),                       //                                                                   .writedata
		.Audio_Subsystem_audio_slave_address                                      (mm_interconnect_0_audio_subsystem_audio_slave_address),          //                                        Audio_Subsystem_audio_slave.address
		.Audio_Subsystem_audio_slave_write                                        (mm_interconnect_0_audio_subsystem_audio_slave_write),            //                                                                   .write
		.Audio_Subsystem_audio_slave_read                                         (mm_interconnect_0_audio_subsystem_audio_slave_read),             //                                                                   .read
		.Audio_Subsystem_audio_slave_readdata                                     (mm_interconnect_0_audio_subsystem_audio_slave_readdata),         //                                                                   .readdata
		.Audio_Subsystem_audio_slave_writedata                                    (mm_interconnect_0_audio_subsystem_audio_slave_writedata),        //                                                                   .writedata
		.Audio_Subsystem_audio_slave_chipselect                                   (mm_interconnect_0_audio_subsystem_audio_slave_chipselect),       //                                                                   .chipselect
		.AV_Config_avalon_av_config_slave_address                                 (mm_interconnect_0_av_config_avalon_av_config_slave_address),     //                                   AV_Config_avalon_av_config_slave.address
		.AV_Config_avalon_av_config_slave_write                                   (mm_interconnect_0_av_config_avalon_av_config_slave_write),       //                                                                   .write
		.AV_Config_avalon_av_config_slave_read                                    (mm_interconnect_0_av_config_avalon_av_config_slave_read),        //                                                                   .read
		.AV_Config_avalon_av_config_slave_readdata                                (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),    //                                                                   .readdata
		.AV_Config_avalon_av_config_slave_writedata                               (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),   //                                                                   .writedata
		.AV_Config_avalon_av_config_slave_byteenable                              (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),  //                                                                   .byteenable
		.AV_Config_avalon_av_config_slave_waitrequest                             (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest), //                                                                   .waitrequest
		.collide_finish_s1_address                                                (mm_interconnect_0_collide_finish_s1_address),                    //                                                  collide_finish_s1.address
		.collide_finish_s1_readdata                                               (mm_interconnect_0_collide_finish_s1_readdata),                   //                                                                   .readdata
		.init_finish_s1_address                                                   (mm_interconnect_0_init_finish_s1_address),                       //                                                     init_finish_s1.address
		.init_finish_s1_readdata                                                  (mm_interconnect_0_init_finish_s1_readdata),                      //                                                                   .readdata
		.init_ship_s1_address                                                     (mm_interconnect_0_init_ship_s1_address),                         //                                                       init_ship_s1.address
		.init_ship_s1_write                                                       (mm_interconnect_0_init_ship_s1_write),                           //                                                                   .write
		.init_ship_s1_readdata                                                    (mm_interconnect_0_init_ship_s1_readdata),                        //                                                                   .readdata
		.init_ship_s1_writedata                                                   (mm_interconnect_0_init_ship_s1_writedata),                       //                                                                   .writedata
		.init_ship_s1_chipselect                                                  (mm_interconnect_0_init_ship_s1_chipselect),                      //                                                                   .chipselect
		.move_trace_finish_s1_address                                             (mm_interconnect_0_move_trace_finish_s1_address),                 //                                               move_trace_finish_s1.address
		.move_trace_finish_s1_readdata                                            (mm_interconnect_0_move_trace_finish_s1_readdata),                //                                                                   .readdata
		.n0_from_hps_s1_address                                                   (mm_interconnect_0_n0_from_hps_s1_address),                       //                                                     n0_from_hps_s1.address
		.n0_from_hps_s1_write                                                     (mm_interconnect_0_n0_from_hps_s1_write),                         //                                                                   .write
		.n0_from_hps_s1_readdata                                                  (mm_interconnect_0_n0_from_hps_s1_readdata),                      //                                                                   .readdata
		.n0_from_hps_s1_writedata                                                 (mm_interconnect_0_n0_from_hps_s1_writedata),                     //                                                                   .writedata
		.n0_from_hps_s1_chipselect                                                (mm_interconnect_0_n0_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.ne_from_hps_s1_address                                                   (mm_interconnect_0_ne_from_hps_s1_address),                       //                                                     ne_from_hps_s1.address
		.ne_from_hps_s1_write                                                     (mm_interconnect_0_ne_from_hps_s1_write),                         //                                                                   .write
		.ne_from_hps_s1_readdata                                                  (mm_interconnect_0_ne_from_hps_s1_readdata),                      //                                                                   .readdata
		.ne_from_hps_s1_writedata                                                 (mm_interconnect_0_ne_from_hps_s1_writedata),                     //                                                                   .writedata
		.ne_from_hps_s1_chipselect                                                (mm_interconnect_0_ne_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.nn_from_hps_s1_address                                                   (mm_interconnect_0_nn_from_hps_s1_address),                       //                                                     nn_from_hps_s1.address
		.nn_from_hps_s1_write                                                     (mm_interconnect_0_nn_from_hps_s1_write),                         //                                                                   .write
		.nn_from_hps_s1_readdata                                                  (mm_interconnect_0_nn_from_hps_s1_readdata),                      //                                                                   .readdata
		.nn_from_hps_s1_writedata                                                 (mm_interconnect_0_nn_from_hps_s1_writedata),                     //                                                                   .writedata
		.nn_from_hps_s1_chipselect                                                (mm_interconnect_0_nn_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.nne_from_hps_s1_address                                                  (mm_interconnect_0_nne_from_hps_s1_address),                      //                                                    nne_from_hps_s1.address
		.nne_from_hps_s1_write                                                    (mm_interconnect_0_nne_from_hps_s1_write),                        //                                                                   .write
		.nne_from_hps_s1_readdata                                                 (mm_interconnect_0_nne_from_hps_s1_readdata),                     //                                                                   .readdata
		.nne_from_hps_s1_writedata                                                (mm_interconnect_0_nne_from_hps_s1_writedata),                    //                                                                   .writedata
		.nne_from_hps_s1_chipselect                                               (mm_interconnect_0_nne_from_hps_s1_chipselect),                   //                                                                   .chipselect
		.nnw_from_hps_s1_address                                                  (mm_interconnect_0_nnw_from_hps_s1_address),                      //                                                    nnw_from_hps_s1.address
		.nnw_from_hps_s1_write                                                    (mm_interconnect_0_nnw_from_hps_s1_write),                        //                                                                   .write
		.nnw_from_hps_s1_readdata                                                 (mm_interconnect_0_nnw_from_hps_s1_readdata),                     //                                                                   .readdata
		.nnw_from_hps_s1_writedata                                                (mm_interconnect_0_nnw_from_hps_s1_writedata),                    //                                                                   .writedata
		.nnw_from_hps_s1_chipselect                                               (mm_interconnect_0_nnw_from_hps_s1_chipselect),                   //                                                                   .chipselect
		.ns_from_hps_s1_address                                                   (mm_interconnect_0_ns_from_hps_s1_address),                       //                                                     ns_from_hps_s1.address
		.ns_from_hps_s1_write                                                     (mm_interconnect_0_ns_from_hps_s1_write),                         //                                                                   .write
		.ns_from_hps_s1_readdata                                                  (mm_interconnect_0_ns_from_hps_s1_readdata),                      //                                                                   .readdata
		.ns_from_hps_s1_writedata                                                 (mm_interconnect_0_ns_from_hps_s1_writedata),                     //                                                                   .writedata
		.ns_from_hps_s1_chipselect                                                (mm_interconnect_0_ns_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.nse_from_hps_s1_address                                                  (mm_interconnect_0_nse_from_hps_s1_address),                      //                                                    nse_from_hps_s1.address
		.nse_from_hps_s1_write                                                    (mm_interconnect_0_nse_from_hps_s1_write),                        //                                                                   .write
		.nse_from_hps_s1_readdata                                                 (mm_interconnect_0_nse_from_hps_s1_readdata),                     //                                                                   .readdata
		.nse_from_hps_s1_writedata                                                (mm_interconnect_0_nse_from_hps_s1_writedata),                    //                                                                   .writedata
		.nse_from_hps_s1_chipselect                                               (mm_interconnect_0_nse_from_hps_s1_chipselect),                   //                                                                   .chipselect
		.nsw_from_hps_s1_address                                                  (mm_interconnect_0_nsw_from_hps_s1_address),                      //                                                    nsw_from_hps_s1.address
		.nsw_from_hps_s1_write                                                    (mm_interconnect_0_nsw_from_hps_s1_write),                        //                                                                   .write
		.nsw_from_hps_s1_readdata                                                 (mm_interconnect_0_nsw_from_hps_s1_readdata),                     //                                                                   .readdata
		.nsw_from_hps_s1_writedata                                                (mm_interconnect_0_nsw_from_hps_s1_writedata),                    //                                                                   .writedata
		.nsw_from_hps_s1_chipselect                                               (mm_interconnect_0_nsw_from_hps_s1_chipselect),                   //                                                                   .chipselect
		.nw_from_hps_s1_address                                                   (mm_interconnect_0_nw_from_hps_s1_address),                       //                                                     nw_from_hps_s1.address
		.nw_from_hps_s1_write                                                     (mm_interconnect_0_nw_from_hps_s1_write),                         //                                                                   .write
		.nw_from_hps_s1_readdata                                                  (mm_interconnect_0_nw_from_hps_s1_readdata),                      //                                                                   .readdata
		.nw_from_hps_s1_writedata                                                 (mm_interconnect_0_nw_from_hps_s1_writedata),                     //                                                                   .writedata
		.nw_from_hps_s1_chipselect                                                (mm_interconnect_0_nw_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.pipes_s1_address                                                         (mm_interconnect_0_pipes_s1_address),                             //                                                           pipes_s1.address
		.pipes_s1_readdata                                                        (mm_interconnect_0_pipes_s1_readdata),                            //                                                                   .readdata
		.print_finish_s1_address                                                  (mm_interconnect_0_print_finish_s1_address),                      //                                                    print_finish_s1.address
		.print_finish_s1_readdata                                                 (mm_interconnect_0_print_finish_s1_readdata),                     //                                                                   .readdata
		.reset_lb_s1_address                                                      (mm_interconnect_0_reset_lb_s1_address),                          //                                                        reset_lb_s1.address
		.reset_lb_s1_write                                                        (mm_interconnect_0_reset_lb_s1_write),                            //                                                                   .write
		.reset_lb_s1_readdata                                                     (mm_interconnect_0_reset_lb_s1_readdata),                         //                                                                   .readdata
		.reset_lb_s1_writedata                                                    (mm_interconnect_0_reset_lb_s1_writedata),                        //                                                                   .writedata
		.reset_lb_s1_chipselect                                                   (mm_interconnect_0_reset_lb_s1_chipselect),                       //                                                                   .chipselect
		.ship_x_s1_address                                                        (mm_interconnect_0_ship_x_s1_address),                            //                                                          ship_x_s1.address
		.ship_x_s1_write                                                          (mm_interconnect_0_ship_x_s1_write),                              //                                                                   .write
		.ship_x_s1_readdata                                                       (mm_interconnect_0_ship_x_s1_readdata),                           //                                                                   .readdata
		.ship_x_s1_writedata                                                      (mm_interconnect_0_ship_x_s1_writedata),                          //                                                                   .writedata
		.ship_x_s1_chipselect                                                     (mm_interconnect_0_ship_x_s1_chipselect),                         //                                                                   .chipselect
		.ship_y_s1_address                                                        (mm_interconnect_0_ship_y_s1_address),                            //                                                          ship_y_s1.address
		.ship_y_s1_write                                                          (mm_interconnect_0_ship_y_s1_write),                              //                                                                   .write
		.ship_y_s1_readdata                                                       (mm_interconnect_0_ship_y_s1_readdata),                           //                                                                   .readdata
		.ship_y_s1_writedata                                                      (mm_interconnect_0_ship_y_s1_writedata),                          //                                                                   .writedata
		.ship_y_s1_chipselect                                                     (mm_interconnect_0_ship_y_s1_chipselect),                         //                                                                   .chipselect
		.speed_color_finish_s1_address                                            (mm_interconnect_0_speed_color_finish_s1_address),                //                                              speed_color_finish_s1.address
		.speed_color_finish_s1_readdata                                           (mm_interconnect_0_speed_color_finish_s1_readdata),               //                                                                   .readdata
		.start_collide_s1_address                                                 (mm_interconnect_0_start_collide_s1_address),                     //                                                   start_collide_s1.address
		.start_collide_s1_write                                                   (mm_interconnect_0_start_collide_s1_write),                       //                                                                   .write
		.start_collide_s1_readdata                                                (mm_interconnect_0_start_collide_s1_readdata),                    //                                                                   .readdata
		.start_collide_s1_writedata                                               (mm_interconnect_0_start_collide_s1_writedata),                   //                                                                   .writedata
		.start_collide_s1_chipselect                                              (mm_interconnect_0_start_collide_s1_chipselect),                  //                                                                   .chipselect
		.start_init_s1_address                                                    (mm_interconnect_0_start_init_s1_address),                        //                                                      start_init_s1.address
		.start_init_s1_write                                                      (mm_interconnect_0_start_init_s1_write),                          //                                                                   .write
		.start_init_s1_readdata                                                   (mm_interconnect_0_start_init_s1_readdata),                       //                                                                   .readdata
		.start_init_s1_writedata                                                  (mm_interconnect_0_start_init_s1_writedata),                      //                                                                   .writedata
		.start_init_s1_chipselect                                                 (mm_interconnect_0_start_init_s1_chipselect),                     //                                                                   .chipselect
		.start_move_trace_s1_address                                              (mm_interconnect_0_start_move_trace_s1_address),                  //                                                start_move_trace_s1.address
		.start_move_trace_s1_write                                                (mm_interconnect_0_start_move_trace_s1_write),                    //                                                                   .write
		.start_move_trace_s1_readdata                                             (mm_interconnect_0_start_move_trace_s1_readdata),                 //                                                                   .readdata
		.start_move_trace_s1_writedata                                            (mm_interconnect_0_start_move_trace_s1_writedata),                //                                                                   .writedata
		.start_move_trace_s1_chipselect                                           (mm_interconnect_0_start_move_trace_s1_chipselect),               //                                                                   .chipselect
		.start_print_s1_address                                                   (mm_interconnect_0_start_print_s1_address),                       //                                                     start_print_s1.address
		.start_print_s1_write                                                     (mm_interconnect_0_start_print_s1_write),                         //                                                                   .write
		.start_print_s1_readdata                                                  (mm_interconnect_0_start_print_s1_readdata),                      //                                                                   .readdata
		.start_print_s1_writedata                                                 (mm_interconnect_0_start_print_s1_writedata),                     //                                                                   .writedata
		.start_print_s1_chipselect                                                (mm_interconnect_0_start_print_s1_chipselect),                    //                                                                   .chipselect
		.start_speed_color_s1_address                                             (mm_interconnect_0_start_speed_color_s1_address),                 //                                               start_speed_color_s1.address
		.start_speed_color_s1_write                                               (mm_interconnect_0_start_speed_color_s1_write),                   //                                                                   .write
		.start_speed_color_s1_readdata                                            (mm_interconnect_0_start_speed_color_s1_readdata),                //                                                                   .readdata
		.start_speed_color_s1_writedata                                           (mm_interconnect_0_start_speed_color_s1_writedata),               //                                                                   .writedata
		.start_speed_color_s1_chipselect                                          (mm_interconnect_0_start_speed_color_s1_chipselect),              //                                                                   .chipselect
		.start_stream_s1_address                                                  (mm_interconnect_0_start_stream_s1_address),                      //                                                    start_stream_s1.address
		.start_stream_s1_write                                                    (mm_interconnect_0_start_stream_s1_write),                        //                                                                   .write
		.start_stream_s1_readdata                                                 (mm_interconnect_0_start_stream_s1_readdata),                     //                                                                   .readdata
		.start_stream_s1_writedata                                                (mm_interconnect_0_start_stream_s1_writedata),                    //                                                                   .writedata
		.start_stream_s1_chipselect                                               (mm_interconnect_0_start_stream_s1_chipselect),                   //                                                                   .chipselect
		.stream_finish_s1_address                                                 (mm_interconnect_0_stream_finish_s1_address),                     //                                                   stream_finish_s1.address
		.stream_finish_s1_readdata                                                (mm_interconnect_0_stream_finish_s1_readdata),                    //                                                                   .readdata
		.test_data_s1_address                                                     (mm_interconnect_0_test_data_s1_address),                         //                                                       test_data_s1.address
		.test_data_s1_write                                                       (mm_interconnect_0_test_data_s1_write),                           //                                                                   .write
		.test_data_s1_readdata                                                    (mm_interconnect_0_test_data_s1_readdata),                        //                                                                   .readdata
		.test_data_s1_writedata                                                   (mm_interconnect_0_test_data_s1_writedata),                       //                                                                   .writedata
		.test_data_s1_chipselect                                                  (mm_interconnect_0_test_data_s1_chipselect),                      //                                                                   .chipselect
		.ux_from_hps_s1_address                                                   (mm_interconnect_0_ux_from_hps_s1_address),                       //                                                     ux_from_hps_s1.address
		.ux_from_hps_s1_write                                                     (mm_interconnect_0_ux_from_hps_s1_write),                         //                                                                   .write
		.ux_from_hps_s1_readdata                                                  (mm_interconnect_0_ux_from_hps_s1_readdata),                      //                                                                   .readdata
		.ux_from_hps_s1_writedata                                                 (mm_interconnect_0_ux_from_hps_s1_writedata),                     //                                                                   .writedata
		.ux_from_hps_s1_chipselect                                                (mm_interconnect_0_ux_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.ux_in_s1_address                                                         (mm_interconnect_0_ux_in_s1_address),                             //                                                           ux_in_s1.address
		.ux_in_s1_readdata                                                        (mm_interconnect_0_ux_in_s1_readdata),                            //                                                                   .readdata
		.uy_from_hps_s1_address                                                   (mm_interconnect_0_uy_from_hps_s1_address),                       //                                                     uy_from_hps_s1.address
		.uy_from_hps_s1_write                                                     (mm_interconnect_0_uy_from_hps_s1_write),                         //                                                                   .write
		.uy_from_hps_s1_readdata                                                  (mm_interconnect_0_uy_from_hps_s1_readdata),                      //                                                                   .readdata
		.uy_from_hps_s1_writedata                                                 (mm_interconnect_0_uy_from_hps_s1_writedata),                     //                                                                   .writedata
		.uy_from_hps_s1_chipselect                                                (mm_interconnect_0_uy_from_hps_s1_chipselect),                    //                                                                   .chipselect
		.uy_in_s1_address                                                         (mm_interconnect_0_uy_in_s1_address),                             //                                                           uy_in_s1.address
		.uy_in_s1_readdata                                                        (mm_interconnect_0_uy_in_s1_readdata),                            //                                                                   .readdata
		.write_address_init_s1_address                                            (mm_interconnect_0_write_address_init_s1_address),                //                                              write_address_init_s1.address
		.write_address_init_s1_write                                              (mm_interconnect_0_write_address_init_s1_write),                  //                                                                   .write
		.write_address_init_s1_readdata                                           (mm_interconnect_0_write_address_init_s1_readdata),               //                                                                   .readdata
		.write_address_init_s1_writedata                                          (mm_interconnect_0_write_address_init_s1_writedata),              //                                                                   .writedata
		.write_address_init_s1_chipselect                                         (mm_interconnect_0_write_address_init_s1_chipselect),             //                                                                   .chipselect
		.x_fish1_s1_address                                                       (mm_interconnect_0_x_fish1_s1_address),                           //                                                         x_fish1_s1.address
		.x_fish1_s1_write                                                         (mm_interconnect_0_x_fish1_s1_write),                             //                                                                   .write
		.x_fish1_s1_readdata                                                      (mm_interconnect_0_x_fish1_s1_readdata),                          //                                                                   .readdata
		.x_fish1_s1_writedata                                                     (mm_interconnect_0_x_fish1_s1_writedata),                         //                                                                   .writedata
		.x_fish1_s1_chipselect                                                    (mm_interconnect_0_x_fish1_s1_chipselect),                        //                                                                   .chipselect
		.x_fish2_s1_address                                                       (mm_interconnect_0_x_fish2_s1_address),                           //                                                         x_fish2_s1.address
		.x_fish2_s1_write                                                         (mm_interconnect_0_x_fish2_s1_write),                             //                                                                   .write
		.x_fish2_s1_readdata                                                      (mm_interconnect_0_x_fish2_s1_readdata),                          //                                                                   .readdata
		.x_fish2_s1_writedata                                                     (mm_interconnect_0_x_fish2_s1_writedata),                         //                                                                   .writedata
		.x_fish2_s1_chipselect                                                    (mm_interconnect_0_x_fish2_s1_chipselect),                        //                                                                   .chipselect
		.y_fish1_s1_address                                                       (mm_interconnect_0_y_fish1_s1_address),                           //                                                         y_fish1_s1.address
		.y_fish1_s1_write                                                         (mm_interconnect_0_y_fish1_s1_write),                             //                                                                   .write
		.y_fish1_s1_readdata                                                      (mm_interconnect_0_y_fish1_s1_readdata),                          //                                                                   .readdata
		.y_fish1_s1_writedata                                                     (mm_interconnect_0_y_fish1_s1_writedata),                         //                                                                   .writedata
		.y_fish1_s1_chipselect                                                    (mm_interconnect_0_y_fish1_s1_chipselect),                        //                                                                   .chipselect
		.y_fish2_s1_address                                                       (mm_interconnect_0_y_fish2_s1_address),                           //                                                         y_fish2_s1.address
		.y_fish2_s1_write                                                         (mm_interconnect_0_y_fish2_s1_write),                             //                                                                   .write
		.y_fish2_s1_readdata                                                      (mm_interconnect_0_y_fish2_s1_readdata),                          //                                                                   .readdata
		.y_fish2_s1_writedata                                                     (mm_interconnect_0_y_fish2_s1_writedata),                         //                                                                   .writedata
		.y_fish2_s1_chipselect                                                    (mm_interconnect_0_y_fish2_s1_chipselect)                         //                                                                   .chipselect
	);

	Computer_System_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (arm_a9_hps_f2h_irq0_irq)   //    sender.irq
	);

	Computer_System_irq_mapper_001 irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),    // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),  // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (system_pll_reset_source_reset),      // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
